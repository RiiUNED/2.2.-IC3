---------------------------------------------------------
-- Entity de Funcion (x, y, z) = (F, G)
library IEEE;
use IEEE.std_logic_1164.all;

entity funcFG is
    port ( F, G: out std_logic; x, y, z: in std_logic);
end entity funcFG;
---------------------------------------------------------
